`timescale 1ns / 1ps

module InstructionDecode(
    input [31:0] instruction,
    output reg [53:0] code
);
    wire [5:0] op;
    wire [5:0] func;
    assign op = instruction[31:26];
    assign func = instruction[5:0];

    always @ *
    begin
        code <= 54'b0;
        casez({op, func})
            12'b000000_100000: code[0]  <= 1'b1; //ADD     0
            12'b000000_100001: code[1]  <= 1'b1; //ADDU    1
            12'b000000_100010: code[2]  <= 1'b1; //SUB     2  
            12'b000000_100011: code[3]  <= 1'b1; //SUBU    3
            12'b000000_100100: code[4]  <= 1'b1; //AND     4
            12'b000000_100101: code[5]  <= 1'b1; //OR      5
            12'b000000_100110: code[6]  <= 1'b1; //XOR     6
            12'b000000_100111: code[7]  <= 1'b1; //NOR     7
            12'b000000_101010: code[8]  <= 1'b1; //SLT     8
            12'b000000_101011: code[9]  <= 1'b1; //SLTU    9
            12'b000000_000000: code[10] <= 1'b1; //SLL     10
            12'b000000_000010: code[11] <= 1'b1; //SRL     11
            12'b000000_000011: code[12] <= 1'b1; //SRA     12
            12'b000000_000100: code[13] <= 1'b1; //SLLV    13
            12'b000000_000110: code[14] <= 1'b1; //SRLV    14
            12'b000000_000111: code[15] <= 1'b1; //SRAV    15
            12'b000000_001000: code[16] <= 1'b1; //JR      16
            12'b001000_??????: code[17] <= 1'b1; //ADDI    17
            12'b001001_??????: code[18] <= 1'b1; //ADDIU   18
            12'b001100_??????: code[19] <= 1'b1; //ANDI    19
            12'b001101_??????: code[20] <= 1'b1; //ORI     20
            12'b001110_??????: code[21] <= 1'b1; //XORI    21
            12'b100011_??????: code[22] <= 1'b1; //LW      22
            12'b101011_??????: code[23] <= 1'b1; //SW      23
            12'b000100_??????: code[24] <= 1'b1; //BEQ     24
            12'b000101_??????: code[25] <= 1'b1; //BNE     25
            12'b001010_??????: code[26] <= 1'b1; //SLTI    26
            12'b001011_??????: code[27] <= 1'b1; //SLTIU   27
            12'b001111_??????: code[28] <= 1'b1; //LUI     28
            12'b000010_??????: code[29] <= 1'b1; //J       29
            12'b000011_??????: code[30] <= 1'b1; //JAL     30
            12'b011100_100000: code[31] <= 1'b1; //CLZ     31
            12'b000000_011011: code[32] <= 1'b1; //DIVU    32
            12'b010000_011000: code[33] <= 1'b1; //ERET    33
            12'b000000_001001: code[34] <= 1'b1; //JALR    34
            12'b100000_??????: code[35] <= 1'b1; //LB      35
            12'b100100_??????: code[36] <= 1'b1; //LBU     36
            12'b100101_??????: code[37] <= 1'b1; //LHU     37
            12'b101000_??????: code[38] <= 1'b1; //SB      38
            12'b101001_??????: code[39] <= 1'b1; //SH      39
            12'b100001_??????: code[40] <= 1'b1; //LH      40
            12'b010000_000000: code[41] <= 1'b1; //MFC0    41*
            12'b000000_010000: code[42] <= 1'b1; //MFHI    42
            12'b000000_010010: code[43] <= 1'b1; //MFLO    43
            12'b010000_000000: code[44] <= 1'b1; //MTC0    44*
            12'b000000_010001: code[45] <= 1'b1; //MTHI    45
            12'b000000_010011: code[46] <= 1'b1; //MTLO    46
            12'b011100_000010: code[47] <= 1'b1; //MUL     47
            12'b000000_011001: code[48] <= 1'b1; //MULTU   48
            12'b000000_001100: code[49] <= 1'b1; //SYSCALL 49
            12'b000000_110100: code[50] <= 1'b1; //TEQ     50
            12'b000001_??????: code[51] <= 1'b1; //BGEZ    51
            12'b000000_001101: code[52] <= 1'b1; //BREAK   52
            12'b000000_011010: code[53] <= 1'b1; //DIV     53
            default:           code <= 54'b0;
        endcase
    end
endmodule
